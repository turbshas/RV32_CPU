`define REG_ADDR_WIDTH 5
`define REGISTER_X0 `REG_ADDR_WIDTH'b0
`define REG_WIDTH 32
